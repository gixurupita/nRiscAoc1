module nRisc (
    ports
);
    
endmodule