module Processador_nRisc (Clock, Reset, RaidaPC, CamposInst, EndMemoria, DadoMemoria);
    input wire
endmodule