module Processador_nRisc (clock, reset, saidaPC, camposInst, endMemoria, dadoMemoria);
    input wire
endmodule